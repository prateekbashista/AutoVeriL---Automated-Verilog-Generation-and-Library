module half_add(input a, input b, output s, output cout); 

assign s = a ^ b;
assign s = a & b;
endmodule